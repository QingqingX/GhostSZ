`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/01/2019 11:42:50 AM
// Design Name: 
// Module Name: fpaddsub
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module aaa(
    input add_sub,
    input clock,
    input [31:0] dataa,
    input [31:0] datab,
    input [31:0] result
    );
endmodule
