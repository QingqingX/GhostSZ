`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/10/2019 04:06:31 PM
// Design Name: 
// Module Name: mux128
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux128(
    input aclr,
	input clock,
	input [31:0] data0x,
	input [31:0] data10x,
	input [31:0] data11x,
	input [31:0] data12x,
	input [31:0] data13x,
    input [31:0] data14x,
	input [31:0] data15x,
	input [31:0] data16x,
	input [31:0] data17x,
	input [31:0] data18x,
	input [31:0] data19x,
	input [31:0] data1x,
	input [31:0] data20x,
	input [31:0] data21x,
	input [31:0] data22x,
	input [31:0] data23x,
	input [31:0] data24x,
	input [31:0] data25x,
	input [31:0] data26x,
	input [31:0] data27x,
	input [31:0] data28x,
	input [31:0] data29x,
	input [31:0] data2x,
	input [31:0] data30x,
	input [31:0] data31x,
	input [31:0] data32x,
	input [31:0] data33x,
	input [31:0] data34x,
	input [31:0] data35x,
	input [31:0] data36x,
	input [31:0] data37x,
	input [31:0] data38x,
	input [31:0] data39x,
	input [31:0] data3x,
	input [31:0] data40x,
	input [31:0] data41x,
	input [31:0] data42x,
	input [31:0] data43x,
	input [31:0] data44x,
	input [31:0] data45x,
	input [31:0] data46x,
	input [31:0] data47x,
	input [31:0] data48x,
	input [31:0] data49x,
	input [31:0] data50x,
    input [31:0] data51x,
    input [31:0] data52x,
    input [31:0] data53x,
    input [31:0] data54x,
    input [31:0] data55x,
    input [31:0] data56x,
    input [31:0] data57x,
    input [31:0] data58x,
    input [31:0] data59x,
    input [31:0] data60x,
    input [31:0] data61x,
    input [31:0] data62x,
    input [31:0] data63x,
	input [31:0] data4x,
	input [31:0] data5x,
	input [31:0] data6x,
	input [31:0] data7x,
	input [31:0] data8x,
	input [31:0] data9x,
		
    input [31:0] data0y,
    input [31:0] data10y,
    input [31:0] data11y,
    input [31:0] data12y,
    input [31:0] data13y,
    input [31:0] data14y,
    input [31:0] data15y,
    input [31:0] data16y,
    input [31:0] data17y,
    input [31:0] data18y,
    input [31:0] data19y,
    input [31:0] data1y,
    input [31:0] data20y,
    input [31:0] data21y,
    input [31:0] data22y,
    input [31:0] data23y,
    input [31:0] data24y,
    input [31:0] data25y,
    input [31:0] data26y,
    input [31:0] data27y,
    input [31:0] data28y,
    input [31:0] data29y,
    input [31:0] data2y,
    input [31:0] data30y,
    input [31:0] data31y,
    input [31:0] data32y,
    input [31:0] data33y,
    input [31:0] data34y,
    input [31:0] data35y,
    input [31:0] data36y,
    input [31:0] data37y,
    input [31:0] data38y,
    input [31:0] data39y,
    input [31:0] data3y,
    input [31:0] data40y,
    input [31:0] data41y,
    input [31:0] data42y,
    input [31:0] data43y,
    input [31:0] data44y,
    input [31:0] data45y,
    input [31:0] data46y,
    input [31:0] data47y,
    input [31:0] data48y,
    input [31:0] data49y,
    input [31:0] data50y,
    input [31:0] data51y,
    input [31:0] data52y,
    input [31:0] data53y,
    input [31:0] data54y,
    input [31:0] data55y,
    input [31:0] data56y,
    input [31:0] data57y,
    input [31:0] data58y,
    input [31:0] data59y,
    input [31:0] data60y,
    input [31:0] data61y,
    input [31:0] data62y,
    input [31:0] data63y,
    input [31:0] data4y,
    input [31:0] data5y,
    input [31:0] data6y,
    input [31:0] data7y,
    input [31:0] data8y,
    input [31:0] data9y,
    
	input [6:0] sel,
	output [31:0] result
    );
    
wire [31:0] result_x, result_y;
mux64  muxx(
        aclr,
        clock,
        data0x,
        data10x,
        data11x,
        data12x,
        data13x,
        data14x,
        data15x,
        data16x,
        data17x,
        data18x,
        data19x,
        data1x,
        data20x,
        data21x,
        data22x,
        data23x,
        data24x,
        data25x,
        data26x,
        data27x,
        data28x,
        data29x,
        data2x,
        data30x,
        data31x,
        data32x,
        data33x,
        data34x,
        data35x,
        data36x,
        data37x,
        data38x,
        data39x,
        data3x,
        data40x,
        data41x,
        data42x,
        data43x,
        data44x,
        data45x,
        data46x,
        data47x,
        data48x,
        data49x,
        data50x,
        data51x,
        data52x,
        data53x,
        data54x,
        data55x,
        data56x,
        data57x,
        data58x,
        data59x,
        data60x,
        data61x,
        data62x,
        data63x,
        data4x,
        data5x,
        data6x,
        data7x,
        data8x,
        data9x,
        sel[5:0],
         result_x
        );    
mux64  muxy(
        aclr,
        clock,
        data0y,
        data10y,
        data11y,
        data12y,
        data13y,
        data14y,
        data15y,
        data16y,
        data17y,
        data18y,
        data19y,
        data1y,
        data20y,
        data21y,
        data22y,
        data23y,
        data24y,
        data25y,
        data26y,
        data27y,
        data28y,
        data29y,
        data2y,
        data30y,
        data31y,
        data32y,
        data33y,
        data34y,
        data35y,
        data36y,
        data37y,
        data38y,
        data39y,
        data3y,
        data40y,
        data41y,
        data42y,
        data43y,
        data44y,
        data45y,
        data46y,
        data47y,
        data48y,
        data49y,
        data50y,
        data51y,
        data52y,
        data53y,
        data54y,
        data55y,
        data56y,
        data57y,
        data58y,
        data59y,
        data60y,
        data61y,
        data62y,
        data63y,
        data4y,
        data5y,
        data6y,
        data7y,
        data8y,
        data9y,
        sel[5:0],
         result_y
        ); 

assign result = sel[6]? result_y: result_x;

endmodule
