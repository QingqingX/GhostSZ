`timescale 1 ns / 100 ps

module sz_inner_tb1;
reg rst;
reg clk;
reg [31:0]  data_in;
wire [1:0] data_out;
wire [31:0] phase3_data_out;
wire [9:0] phase2_data_out;
wire phase2_valid, phase3_valid;

sz_inner sz0(
    rst,
    clk,
    data_in,
	data_out,
	phase2_data_out,
	phase2_valid,
	phase3_data_out,
	phase3_valid
);


always #1 clk=~clk;

//integer               data_file    ; // file handler
//integer               scan_file    ; // file handler
//reg [31:0] captured_data;

//integer f;

initial begin
	//f = $fopen("output.txt","w");
  //data_file = $fopen("/home/qx/compress/in.txt", "r");
  //if (data_file == 0) begin
  //  $display("data_file handle was NULL");
  //  $finish;
  //end
  
  clk=0;
  rst=1;
#11 rst=0;
 data_in=32'h3e702c81;
#2 data_in=32'h3e702625;
#2 data_in=32'h3e7022c4;
#2 data_in=32'h3e702322;
#2 data_in=32'h3e702491;
#2 data_in=32'h3e702a25;
#2 data_in=32'h3e703406;
#2 data_in=32'h3e7038db;
#2 data_in=32'h3e702c81;
#2 data_in=32'h3e702625;
#2 data_in=32'h3e7022c4;
#2 data_in=32'h3e702322;
#2 data_in=32'h3e702491;
#2 data_in=32'h3e702a25;
#2 data_in=32'h3e703406;
#2 data_in=32'h3e7038db;
#2 data_in=32'h3e702c81;
#2 data_in=32'h3e702625;
#2 data_in=32'h3e7022c4;
#2 data_in=32'h3e702322;
#2 data_in=32'h3e702491;
#2 data_in=32'h3e702a25;
#2 data_in=32'h3e703406;
#2 data_in=32'h3e7038db;
#2 data_in=32'h3e702c81;
#2 data_in=32'h3e702625;
#2 data_in=32'h3e7022c4;
#2 data_in=32'h3e702322;
#2 data_in=32'h3e702491;
#2 data_in=32'h3e702a25;
#2 data_in=32'h3e703406;
#2 data_in=32'h3e7038db;
#2 data_in=32'h3e702c81;
#2 data_in=32'h3e702625;
#2 data_in=32'h3e7022c4;
#2 data_in=32'h3e702322;
#2 data_in=32'h3e702491;
#2 data_in=32'h3e702a25;
#2 data_in=32'h3e703406;
#2 data_in=32'h3e7038db;
#2 data_in=32'h3e702c81;
#2 data_in=32'h3e702625;
#2 data_in=32'h3e7022c4;
#2 data_in=32'h3e702322;
#2 data_in=32'h3e702491;
#2 data_in=32'h3e702a25;
#2 data_in=32'h3e703406;
#2 data_in=32'h3e7038db;
#2 data_in=32'h3e702c81;
#2 data_in=32'h3e702625;
#2 data_in=32'h3e7022c4;
#2 data_in=32'h3e702322;
#2 data_in=32'h3e702491;
#2 data_in=32'h3e702a25;
#2 data_in=32'h3e703406;
#2 data_in=32'h3e7038db;
#2 data_in=32'h3e702c81;
#2 data_in=32'h3e702625;
#2 data_in=32'h3e7022c4;
#2 data_in=32'h3e702322;
#2 data_in=32'h3e702491;
#2 data_in=32'h3e702a25;
#2 data_in=32'h3e703406;
#2 data_in=32'h3e7038db;
#2 data_in=32'h3e702fa1;
#2 data_in=32'h3e70185e;
#2 data_in=32'h3e6ff733;
#2 data_in=32'h3e6fda19;
#2 data_in=32'h3e6fc8ae;
#2 data_in=32'h3e6fc19a;
#2 data_in=32'h3e6fbf4e;
#2 data_in=32'h3e6fb840;
#2 data_in=32'h3e702fa1;
#2 data_in=32'h3e70185e;
#2 data_in=32'h3e6ff733;
#2 data_in=32'h3e6fda19;
#2 data_in=32'h3e6fc8ae;
#2 data_in=32'h3e6fc19a;
#2 data_in=32'h3e6fbf4e;
#2 data_in=32'h3e6fb840;
#2 data_in=32'h3e702fa1;
#2 data_in=32'h3e70185e;
#2 data_in=32'h3e6ff733;
#2 data_in=32'h3e6fda19;
#2 data_in=32'h3e6fc8ae;
#2 data_in=32'h3e6fc19a;
#2 data_in=32'h3e6fbf4e;
#2 data_in=32'h3e6fb840;
#2 data_in=32'h3e702fa1;
#2 data_in=32'h3e70185e;
#2 data_in=32'h3e6ff733;
#2 data_in=32'h3e6fda19;
#2 data_in=32'h3e6fc8ae;
#2 data_in=32'h3e6fc19a;
#2 data_in=32'h3e6fbf4e;
#2 data_in=32'h3e6fb840;
#2 data_in=32'h3e702fa1;
#2 data_in=32'h3e70185e;
#2 data_in=32'h3e6ff733;
#2 data_in=32'h3e6fda19;
#2 data_in=32'h3e6fc8ae;
#2 data_in=32'h3e6fc19a;
#2 data_in=32'h3e6fbf4e;
#2 data_in=32'h3e6fb840;
#2 data_in=32'h3e702fa1;
#2 data_in=32'h3e70185e;
#2 data_in=32'h3e6ff733;
#2 data_in=32'h3e6fda19;
#2 data_in=32'h3e6fc8ae;
#2 data_in=32'h3e6fc19a;
#2 data_in=32'h3e6fbf4e;
#2 data_in=32'h3e6fb840;
#2 data_in=32'h3e702fa1;
#2 data_in=32'h3e70185e;
#2 data_in=32'h3e6ff733;
#2 data_in=32'h3e6fda19;
#2 data_in=32'h3e6fc8ae;
#2 data_in=32'h3e6fc19a;
#2 data_in=32'h3e6fbf4e;
#2 data_in=32'h3e6fb840;
#2 data_in=32'h3e702fa1;
#2 data_in=32'h3e70185e;
#2 data_in=32'h3e6ff733;
#2 data_in=32'h3e6fda19;
#2 data_in=32'h3e6fc8ae;
#2 data_in=32'h3e6fc19a;
#2 data_in=32'h3e6fbf4e;
#2 data_in=32'h3e6fb840;
#2 data_in=32'h3e6fa227;
#2 data_in=32'h3e6f70b9;
#2 data_in=32'h3e6f2b31;
#2 data_in=32'h3e6ee652;
#2 data_in=32'h3e6ea786;
#2 data_in=32'h3e6e777d;
#2 data_in=32'h3e6e4a5b;
#2 data_in=32'h3e6e1228;
#2 data_in=32'h3e6fa227;
#2 data_in=32'h3e6f70b9;
#2 data_in=32'h3e6f2b31;
#2 data_in=32'h3e6ee652;
#2 data_in=32'h3e6ea786;
#2 data_in=32'h3e6e777d;
#2 data_in=32'h3e6e4a5b;
#2 data_in=32'h3e6e1228;
#2 data_in=32'h3e6fa227;
#2 data_in=32'h3e6f70b9;
#2 data_in=32'h3e6f2b31;
#2 data_in=32'h3e6ee652;
#2 data_in=32'h3e6ea786;
#2 data_in=32'h3e6e777d;
#2 data_in=32'h3e6e4a5b;
#2 data_in=32'h3e6e1228;
#2 data_in=32'h3e6fa227;
#2 data_in=32'h3e6f70b9;
#2 data_in=32'h3e6f2b31;
#2 data_in=32'h3e6ee652;
#2 data_in=32'h3e6ea786;
#2 data_in=32'h3e6e777d;
#2 data_in=32'h3e6e4a5b;
#2 data_in=32'h3e6e1228;
#2 data_in=32'h3e6fa227;
#2 data_in=32'h3e6f70b9;
#2 data_in=32'h3e6f2b31;
#2 data_in=32'h3e6ee652;
#2 data_in=32'h3e6ea786;
#2 data_in=32'h3e6e777d;
#2 data_in=32'h3e6e4a5b;
#2 data_in=32'h3e6e1228;
#2 data_in=32'h3e6fa227;
#2 data_in=32'h3e6f70b9;
#2 data_in=32'h3e6f2b31;
#2 data_in=32'h3e6ee652;
#2 data_in=32'h3e6ea786;
#2 data_in=32'h3e6e777d;
#2 data_in=32'h3e6e4a5b;
#2 data_in=32'h3e6e1228;
#2 data_in=32'h3e6fa227;
#2 data_in=32'h3e6f70b9;
#2 data_in=32'h3e6f2b31;
#2 data_in=32'h3e6ee652;
#2 data_in=32'h3e6ea786;
#2 data_in=32'h3e6e777d;
#2 data_in=32'h3e6e4a5b;
#2 data_in=32'h3e6e1228;
#2 data_in=32'h3e6fa227;
#2 data_in=32'h3e6f70b9;
#2 data_in=32'h3e6f2b31;
#2 data_in=32'h3e6ee652;
#2 data_in=32'h3e6ea786;
#2 data_in=32'h3e6e777d;
#2 data_in=32'h3e6e4a5b;
#2 data_in=32'h3e6e1228;
#2 data_in=32'h3e6dca87;
#2 data_in=32'h3e6d723e;
#2 data_in=32'h3e6cf496;
#2 data_in=32'h3e6c3f87;
#2 data_in=32'h3e6b610e;
#2 data_in=32'h3e6a721e;
#2 data_in=32'h3e6972f5;
#2 data_in=32'h3e68784b;
#2 data_in=32'h3e6dca87;
#2 data_in=32'h3e6d723e;
#2 data_in=32'h3e6cf496;
#2 data_in=32'h3e6c3f87;
#2 data_in=32'h3e6b610e;
#2 data_in=32'h3e6a721e;
#2 data_in=32'h3e6972f5;
#2 data_in=32'h3e68784b;
#2 data_in=32'h3e6dca87;
#2 data_in=32'h3e6d723e;
#2 data_in=32'h3e6cf496;
#2 data_in=32'h3e6c3f87;
#2 data_in=32'h3e6b610e;
#2 data_in=32'h3e6a721e;
#2 data_in=32'h3e6972f5;
#2 data_in=32'h3e68784b;
#2 data_in=32'h3e6dca87;
#2 data_in=32'h3e6d723e;
#2 data_in=32'h3e6cf496;
#2 data_in=32'h3e6c3f87;
#2 data_in=32'h3e6b610e;
#2 data_in=32'h3e6a721e;
#2 data_in=32'h3e6972f5;
#2 data_in=32'h3e68784b;
#2 data_in=32'h3e6dca87;
#2 data_in=32'h3e6d723e;
#2 data_in=32'h3e6cf496;
#2 data_in=32'h3e6c3f87;
#2 data_in=32'h3e6b610e;
#2 data_in=32'h3e6a721e;
#2 data_in=32'h3e6972f5;
#2 data_in=32'h3e68784b;
#2 data_in=32'h3e6dca87;
#2 data_in=32'h3e6d723e;
#2 data_in=32'h3e6cf496;
#2 data_in=32'h3e6c3f87;
#2 data_in=32'h3e6b610e;
#2 data_in=32'h3e6a721e;
#2 data_in=32'h3e6972f5;
#2 data_in=32'h3e68784b;
#2 data_in=32'h3e6dca87;
#2 data_in=32'h3e6d723e;
#2 data_in=32'h3e6cf496;
#2 data_in=32'h3e6c3f87;
#2 data_in=32'h3e6b610e;
#2 data_in=32'h3e6a721e;
#2 data_in=32'h3e6972f5;
#2 data_in=32'h3e68784b;
#2 data_in=32'h3e6dca87;
#2 data_in=32'h3e6d723e;
//$fwrite(f,"%b\n",   data_out);
#600 rst=1;
#20 $stop;
end
endmodule
